module ksa16(
    input  [15:0] a,
    input  [15:0] b,
    output [16:0] sum
);
    wire [15:0] g, p;  // generate and propagate
    wire [15:0] c;     // carry signals

    // Generate and Propagate signals
    assign g = a & b;
    assign p = a ^ b;

    // Carry computation (fully expanded)
    assign c[0]  = g[0];
    assign c[1]  = g[1] | (p[1] & g[0]);
    assign c[2]  = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]);
    assign c[3]  = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]);
    assign c[4]  = g[4] | (p[4] & g[3]) | (p[4] & p[3] & g[2]) | (p[4] & p[3] & p[2] & g[1]) | (p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[5]  = g[5] | (p[5] & g[4]) | (p[5] & p[4] & g[3]) | (p[5] & p[4] & p[3] & g[2]) | (p[5] & p[4] & p[3] & p[2] & g[1]) | (p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[6]  = g[6] | (p[6] & g[5]) | (p[6] & p[5] & g[4]) | (p[6] & p[5] & p[4] & g[3]) | (p[6] & p[5] & p[4] & p[3] & g[2]) | (p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[7]  = g[7] | (p[7] & g[6]) | (p[7] & p[6] & g[5]) | (p[7] & p[6] & p[5] & g[4]) | (p[7] & p[6] & p[5] & p[4] & g[3]) | (p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[8]  = g[8] | (p[8] & g[7]) | (p[8] & p[7] & g[6]) | (p[8] & p[7] & p[6] & g[5]) | (p[8] & p[7] & p[6] & p[5] & g[4]) | (p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[9]  = g[9] | (p[9] & g[8]) | (p[9] & p[8] & g[7]) | (p[9] & p[8] & p[7] & g[6]) | (p[9] & p[8] & p[7] & p[6] & g[5]) | (p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[10] = g[10] | (p[10] & g[9]) | (p[10] & p[9] & g[8]) | (p[10] & p[9] & p[8] & g[7]) | (p[10] & p[9] & p[8] & p[7] & g[6]) | (p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[11] = g[11] | (p[11] & g[10]) | (p[11] & p[10] & g[9]) | (p[11] & p[10] & p[9] & g[8]) | (p[11] & p[10] & p[9] & p[8] & g[7]) | (p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]);
    assign c[12] = g[12] | (p[12]&g[11]) | (p[12]&p[11]&g[10]) | (p[12]&p[11]&p[10]&g[9]) | (p[12]&p[11]&p[10]&p[9]&g[8]) | (p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]);
    assign c[13] = g[13] | (p[13]&g[12]) | (p[13]&p[12]&g[11]) | (p[13]&p[12]&p[11]&g[10]) | (p[13]&p[12]&p[11]&p[10]&g[9]) | (p[13]&p[12]&p[11]&p[10]&p[9]&g[8]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]);
    assign c[14] = g[14] | (p[14]&g[13]) | (p[14]&p[13]&g[12]) | (p[14]&p[13]&p[12]&g[11]) | (p[14]&p[13]&p[12]&p[11]&g[10]) | (p[14]&p[13]&p[12]&p[11]&p[10]&g[9]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]);
    assign c[15] = g[15] | (p[15]&g[14]) | (p[15]&p[14]&g[13]) | (p[15]&p[14]&p[13]&g[12]) | (p[15]&p[14]&p[13]&p[12]&g[11]) | (p[15]&p[14]&p[13]&p[12]&p[11]&g[10]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1]) | (p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0]);

    // Final sum computation
    assign sum[0]  = p[0];
    assign sum[1]  = p[1]  ^ c[0];
    assign sum[2]  = p[2]  ^ c[1];
    assign sum[3]  = p[3]  ^ c[2];
    assign sum[4]  = p[4]  ^ c[3];
    assign sum[5]  = p[5]  ^ c[4];
    assign sum[6]  = p[6]  ^ c[5];
    assign sum[7]  = p[7]  ^ c[6];
    assign sum[8]  = p[8]  ^ c[7];
    assign sum[9]  = p[9]  ^ c[8];
    assign sum[10] = p[10] ^ c[9];
    assign sum[11] = p[11] ^ c[10];
    assign sum[12] = p[12] ^ c[11];
    assign sum[13] = p[13] ^ c[12];
    assign sum[14] = p[14] ^ c[13];
    assign sum[15] = p[15] ^ c[14];
    assign sum[16] = c[15];  // final carry-out
endmodule
